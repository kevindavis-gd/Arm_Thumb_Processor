library verilog;
use verilog.vl_types.all;
entity Logic_vlg_vec_tst is
end Logic_vlg_vec_tst;
